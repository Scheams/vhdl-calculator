library ieee;
use ieee.std_logic_1164.all;

architecture rtl of alu is

begin

end rtl;
