library ieee;
use ieee.std_logic_1164.all;

entity tb_alu is
end tb_alu;

architecture sim of tb_alu is

begin

end sim;
